
`timescale 10ns/10ns 

module nop();

endmodule
