
module reg_data_types();

reg scal;
reg [7:0] vect;
reg [7:0] mem [31:0];
integer i;
integer i_mem [7:0];
time t;
time t_mem [3:0];
real r;
realtime rt1, rt2;

endmodule
