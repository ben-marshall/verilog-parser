
module test;
reg [7:0] mema[0:255];
reg arrayb[7:0][0:255];
wire w_array[7:0][5:0];
integer inta[1:64];
time chng_hist[1:1000];
integer t_index;
endmodule
